module GrayScale (
    input [7:0] r,    // 红色分量（0到255）
    input [7:0] g,    // 绿色分量（0到255）
    input [7:0] b,    // 蓝色分量（0到255）
    output reg [7:0] Gray,// 输出灰度值（0到255）
    output  reg [15:0] Gray_1   // 输出变换后的灰度值，16位，以提供更大的范围

//    output reg [15:0] GAO_data // 假设用16位存储灰度值，GAO数据存储
);

// 计算灰度值
always @ (r or g or b) begin
    Gray = (77 * r + 150 * g + 29 * b)>>8; // 使用加权平均法计算灰度
end

// 假设在某个时刻需要存储灰度值到GAO文件中
//always @ (Gray) begin
//    GAO_data = {8'b0, Gray};  // 将8位灰度值存储到16位变量中
//end


    // 常数c，用于调整对数变换的幅度
    parameter c = 256; // 假设c为256，这个值可以根据需要进行调整

    // 查找表，用于近似对数函数
    // 这里只给出了一个简化的示例，实际使用时需要生成更精确的查找表
//    reg [15:0] lut[255:0] = {
//16'd0, 16'd177, 16'd281, 16'd355, 16'd412, 16'd459, 16'd498, 16'd532, 
//16'd562, 16'd589, 16'd614, 16'd636, 16'd657, 16'd676, 16'd693, 16'd710, 
//16'd725, 16'd740, 16'd754, 16'd767, 16'd779, 16'd791, 16'd803, 16'd814, 
//16'd824, 16'd834, 16'd844, 16'd853, 16'd862, 16'd871, 16'd879, 16'd887, 
//16'd895, 16'd903, 16'd910, 16'd917, 16'd924, 16'd931, 16'd938, 16'd944, 
//16'd951, 16'd957, 16'd963, 16'd969, 16'd975, 16'd980, 16'd986, 16'd991, 
//16'd996, 16'd1001, 16'd1007, 16'd1012, 16'd1016, 16'd1021, 16'd1026, 16'd1030, 
//16'd1035, 16'd1039, 16'd1044, 16'd1048, 16'd1052, 16'd1057, 16'd1061, 16'd1065, 
//16'd1069, 16'd1073, 16'd1076, 16'd1080, 16'd1084, 16'd1088, 16'd1091, 16'd1095, 
//16'd1098, 16'd1102, 16'd1105, 16'd1109, 16'd1112, 16'd1115, 16'd1119, 16'd1122, 
//16'd1125, 16'd1128, 16'd1131, 16'd1134, 16'd1137, 16'd1140, 16'd1143, 16'd1146, 
//16'd1149, 16'd1152, 16'd1155, 16'd1158, 16'd1160, 16'd1163, 16'd1166, 16'd1168, 
//16'd1171, 16'd1174, 16'd1176, 16'd1179, 16'd1181, 16'd1184, 16'd1186, 16'd1189, 
//16'd1191, 16'd1194, 16'd1196, 16'd1199, 16'd1201, 16'd1203, 16'd1206, 16'd1208, 
//16'd1210, 16'd1212, 16'd1215, 16'd1217, 16'd1219, 16'd1221, 16'd1223, 16'd1226, 
//16'd1228, 16'd1230, 16'd1232, 16'd1234, 16'd1236, 16'd1238, 16'd1240, 16'd1242, 
//16'd1244, 16'd1246, 16'd1248, 16'd1250, 16'd1252, 16'd1254, 16'd1256, 16'd1258, 
//16'd1260, 16'd1261, 16'd1263, 16'd1265, 16'd1267, 16'd1269, 16'd1270, 16'd1272, 
//16'd1274, 16'd1276, 16'd1278, 16'd1279, 16'd1281, 16'd1283, 16'd1284, 16'd1286, 
//16'd1288, 16'd1289, 16'd1291, 16'd1293, 16'd1294, 16'd1296, 16'd1298, 16'd1299, 
//16'd1301, 16'd1302, 16'd1304, 16'd1306, 16'd1307, 16'd1309, 16'd1310, 16'd1312, 
//16'd1313, 16'd1315, 16'd1316, 16'd1318, 16'd1319, 16'd1321, 16'd1322, 16'd1324, 
//16'd1325, 16'd1327, 16'd1328, 16'd1329, 16'd1331, 16'd1332, 16'd1334, 16'd1335, 
//16'd1336, 16'd1338, 16'd1339, 16'd1341, 16'd1342, 16'd1343, 16'd1345, 16'd1346, 
//16'd1347, 16'd1349, 16'd1350, 16'd1351, 16'd1353, 16'd1354, 16'd1355, 16'd1356, 
//16'd1358, 16'd1359, 16'd1360, 16'd1361, 16'd1363, 16'd1364, 16'd1365, 16'd1366, 
//16'd1368, 16'd1369, 16'd1370, 16'd1371, 16'd1372, 16'd1374, 16'd1375, 16'd1376, 
//16'd1377, 16'd1378, 16'd1380, 16'd1381, 16'd1382, 16'd1383, 16'd1384, 16'd1385, 
//16'd1387, 16'd1388, 16'd1389, 16'd1390, 16'd1391, 16'd1392, 16'd1393, 16'd1394, 
//16'd1395, 16'd1397, 16'd1398, 16'd1399, 16'd1400, 16'd1401, 16'd1402, 16'd1403, 
//16'd1404, 16'd1405, 16'd1406, 16'd1407, 16'd1408, 16'd1409, 16'd1410, 16'd1411, 
//16'd1412, 16'd1413, 16'd1415, 16'd1416, 16'd1417, 16'd1418, 16'd1419, 16'd1420 


//    };

    // 使用查找表进行变换
always @ (Gray) begin
     Gray_1 =  Gray*c ; // 使用加权平均法计算灰度
end
     // 注意：这里实际上没有直接乘以c，因为lut已经包含了c的影响
                                     // 如果要单独调整c，需要修改查找表的生成方式

    // 注意：上面的代码有一个问题，即直接乘以c可能会导致溢出。
    // 在实际实现中，你可能需要对查找表的值进行缩放，或者对结果进行截断/舍入。
    // 此外，由于我们使用了16位输出，因此查找表的值应该被相应地缩放以匹配这个范围。

    // 更精确的实现可能需要使用多个查找表条目来逼近对数函数的不同部分，
    // 或者使用分段线性逼近等方法。

    // 这里的代码主要是为了演示目的，并不是一个精确的对数变换实现。

endmodule

    
//module top(
//    input clk,       // 时钟信号
//    input reset,     // 复位信号
//    input [7:0] r_R_0_in,
//    input [7:0] r_G_0_in,
//    input [7:0] r_B_0_in,
//    output [7:0] Gray_out,
//    output [7:0] r_R_0_out,
//    output [7:0] r_G_0_out,
//    output [7:0] r_B_0_out
//);
 
    // 实例化rgb_to_gray模块


